module {{ module_name }}();

// some code to generate clock


//  --------------------input/output data types-----------

{{ wire_defs }}

//  --------------------module instancces-----------------

{{instances}}

//  --------------------module assignments-----------------

{{ assignments }}

endmodule
